module main 

import memory_hog
import cpu_exhaust 

fn main()  {
	// memory_hog.run()
	// cpu_exhaust.run()
}