module main 

import uuid

fn main()  {
	println(uuid.new())
	println(uuid.new_upper())
}