module cpu_exhaust

pub fn run() {
	go exhaust_single()
	go exhaust_single()
	go exhaust_single()
	go exhaust_single()

	for true {

	}
}

fn exhaust_single() {
	for true {
		
	}
}